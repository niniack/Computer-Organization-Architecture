`include "half-adder.v"

module half_adder_tb;

  reg a = 0;
  reg b = 0;
  wire sum;
  wire carry;

  half_adder ha(
    .a(a),
    .b(b),
    .sum(sum),
    .carry(carry)
  );

  initial begin
    $dumpfile("half-adder.vcd");
    $dumpvars(0, half_adder_tb);

    a = 1'b0;
    b = 1'b0;
    #10;
    a = 1'b0;
    b = 1'b1;
    #10;
    a = 1'b1;
    b = 1'b0;
    #10;
    a = 1'b1;
    b = 1'b1;
    #10;
  end

endmodule
